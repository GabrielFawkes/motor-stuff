library verilog;
use verilog.vl_types.all;
entity test297_vlg_check_tst is
    port(
        slow_clk        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end test297_vlg_check_tst;
