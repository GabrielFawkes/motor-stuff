library verilog;
use verilog.vl_types.all;
entity L297_vlg_check_tst is
    port(
        clk_out         : in     vl_logic;
        control         : in     vl_logic;
        enable          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end L297_vlg_check_tst;
