library verilog;
use verilog.vl_types.all;
entity L297_vlg_vec_tst is
end L297_vlg_vec_tst;
