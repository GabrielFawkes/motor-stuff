library verilog;
use verilog.vl_types.all;
entity test297_vlg_vec_tst is
end test297_vlg_vec_tst;
