library verilog;
use verilog.vl_types.all;
entity test297 is
    port(
        clk             : in     vl_logic;
        slow_clk        : out    vl_logic
    );
end test297;
