library verilog;
use verilog.vl_types.all;
entity L297 is
    port(
        clk             : in     vl_logic;
        restn_in        : in     vl_logic;
        enable          : out    vl_logic;
        clk_out         : out    vl_logic;
        control         : out    vl_logic
    );
end L297;
