library verilog;
use verilog.vl_types.all;
entity L297_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        restn_in        : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end L297_vlg_sample_tst;
